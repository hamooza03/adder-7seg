module hex_7seg_decoder();


