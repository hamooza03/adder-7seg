module tb_hex_7seg_decoder();