module adder_nbit_top();


